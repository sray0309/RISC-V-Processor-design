
`timescale 1ns / 1ps

`define ZERO_WORD  64'h00000000_00000000   
`define REG_BUS    63 : 0     
`define DATA_WIDTH 64
`define INST_ADD   8'h11
